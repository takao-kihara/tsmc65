//`include "POLYPHASE_PATH4_ADC_TEG.v"
//`include "POLYPHASE_PATH4X2_ADC_TEG.v"

module CIC_FILTER_4X2P_ADC_TEG (IN, CLK, CLK_2, CLK_4, RES, ENABLE, OUT);

	parameter BW = 6;

	input CLK, CLK_2, CLK_4, ENABLE, RES;
       input signed [BW-1:0] IN;
	output signed [BW+3:0]OUT;
	wire signed [BW-1:0] OUT01, OUT02, OUT03, OUT04;

	POLYPHASE_PATH4_ADC_TEG POLYPHASE_01(CLK, CLK_2, CLK_4, RES, ENABLE, IN, OUT01, OUT02, OUT03, OUT04);

	POLYPHASE_PATH4X2_ADC_TEG POLYPASE_02(CLK_4, RES, OUT01, OUT02, OUT03, OUT04, OUT);
	
endmodule
